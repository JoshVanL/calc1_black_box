library verilog;
use verilog.vl_types.all;
entity calc1_testbench is
end calc1_testbench;
