library verilog;
use verilog.vl_types.all;
entity test_calc1_tb is
end test_calc1_tb;
