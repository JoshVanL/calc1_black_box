library verilog;
use verilog.vl_types.all;
entity checkers is
end checkers;
