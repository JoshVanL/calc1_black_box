library verilog;
use verilog.vl_types.all;
entity sub_calc1_tb is
end sub_calc1_tb;
